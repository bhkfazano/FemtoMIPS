library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity cache_instrucoes is
	port( end1: in std_logic_vector(31 downto 0);
		clkC: in std_logic;
		dout: out std_logic_vector(31 downto 0));
end cache_instrucoes;

architecture arch_cache_instrucoes of cache_instrucoes is
	type data is array(0 to 65535) of std_logic_vector(7 downto 0);
	
	signal data_mem: data := 
			--(0 => "00100000") & (1 => "00000001") & (2 => "00000000") & (3 => "00001010") & --addi $0, $1, 10
			
			--(4 => "00100000") & (5 => "00100010") & (6 => "00000000") & (7 => "00001011") & --addi $1, $2, 11
			
			--(8 => "00000000") & (9 => "00000000") & (10 => "00000000") & (11 => "00000000") & 
			
			--(12 => "10101100") & (13 => "00000010") & (14 => "00000000") & (15 => "00010000") & --sw $2, 16($0)
			
			--(16 => "10001100") & (17 => "00000110") & (18 => "00000000") & (19 => "00010000") & --lw $6, 16($0)
			
			--(20 => "10101100") & (21 => "00000110") & (22 => "00000000") & (23 => "00000000") & --sw $6, 0($0)
			
			--(4 => "10101100") & (5 => "00000001") & (6 => "00000000") & (7 => "00010000") & --sw $1, 16($0)
			
			--(8 => "10001100") & (9 => "00000110") & (10 => "00000000") & (11 => "00010000") & --lw $6, 16($0)
			
			--(12 => "10101100") & (13 => "00000110") & (14 => "00000000") & (15 => "00000000") & --sw $6, 0($0)
			
			--(24 to 65535 => "00000000");
			
			
			(0 => "00100000") & (1 => "00000001") & (2 => "00000000") & (3 => "00001010") & --addi $0, $1, 10
			
			(4 => "00100000") & (5 => "01100010") & (6 => "00000000") & (7 => "00100000") & --addi $3, $2, 32
			
			--(8 => "00000000") & (9 => "01000000") & (10 => "00000000") & (11 => "00001000") & --jr $2
			--(8 => "00001100") & (9 => "00000000") & (10 => "00000000") & (11 => "00000110") & --jal 24
			--(8 => "00001000") & (9 => "00000000") & (10 => "00000000") & (11 => "00000110") & --j 24
			(8 => "00000000") & (9 => "00000000") & (10 => "00000000") & (11 => "00000000") & 
			
			(12 => "00000000") & (13 => "00000010") & (14 => "00001000") & (15 => "10000000") & --sll $2, $1, 2
			
			(16 => "00000000") & (17 => "00100010") & (18 => "00011000") & (19 => "00100001") & --addu $1, $2, $3
			
			(20 => "00101000") & (21 => "00100100") & (22 => "00000000") & (23 => "10000000") & --slti $1, $4, 128
			
			(24 => "00000000") & (25 => "10000001") & (26 => "00101000") & (27 => "00101010") & --slt $4, $1, $5
			
			(28 => "10101100") & (29 => "00000011") & (30 => "00000000") & (31 => "00010000") & --sw $3, 16($0)
			
			(32 => "10001100") & (33 => "00000110") & (34 => "00000000") & (35 => "00010000") & --lw $6, 16($0)
			
			(36 => "10101100") & (37 => "00000110") & (38 => "00000000") & (39 => "00000000") & --sw $6, 0($0)
			
			(40 => "10001100") & (41 => "00000111") & (42 => "00000000") & (43 => "00000000") & --lw $7, 0($0)
			
			--(44 => "00010100") & (45 => "11000111") & (46 => "00000000") & (47 => "00000001") & --bne $6, $7, 1
			--(44 => "00000000") & (45 => "00000000") & (46 => "00000000") & (47 => "00000000") & 
			(44 => "00100000") & (45 => "11101000") & (46 => "00000000") & (47 => "00000111") & --addi $7, $8, 7
			
			(48 => "00100001") & (49 => "00001000") & (50 => "00000000") & (51 => "00000111") & --addi $8, $8, 7
			
			(52 => "10101100") & (53 => "00001000") & (54 => "00000000") & (55 => "00100000") & --sw $8, 32($0)
			
			(56 to 65535 => "00000000");
			
			--(28 => "10101100") & (29 => "00000101") & (30 => "00000000") & (31 => "00010000") & --sw $5, 16($0)
			
			--(32 => "10001100") & (33 => "00000110") & (34 => "00000000") & (35 => "00010000") & --lw $6, 16($0)
			
			--(36 => "10101100") & (37 => "00000110") & (38 => "00000000") & (39 => "00100000") & --sw $6, 32($0)
			
			--(40 => "10001100") & (41 => "00000111") & (42 => "00000000") & (43 => "00100000") & --lw $7, 32($0)
			
			--(44 => "00100000") & (45 => "11101000") & (46 => "00000000") & (47 => "00000111") & --addi $7, $8, 7
			
			--(48 => "10101100") & (49 => "00001000") & (50 => "00000000") & (51 => "00000000") & --sw $8, 0($0)
			
			--(52 => "00000000") & (53 => "00000000") & (54 => "00000000") & (55 => "00000000") & 
			--(56 => "00000000") & (57 => "00000000") & (58 => "00000000") & (59 => "00000000") & 
			
			--(60 => "10101100") & (61 => "00000001") & (62 => "00000000") & (63 => "00000000") & 
			
			--(8 => "00010000") & (9 => "00100010") & (10 => "00000000") & (11 => "00000001") & --beq $1, $2, 1
			--(16 => "00001100") & (17 => "00000000") & (18 => "00000000") & (19 => "00011100") & --$31 = 20; go to 28
			
			--(others => (others => '0'));
	
	signal sig_dout: std_logic_vector(31 downto 0) := (others => '0');
	
begin
	process is
	begin
		wait until rising_edge (clkC);
		wait for 0.1 ns;
		if (to_integer(unsigned(end1)) < 65536) then
			wait for 4.9 ns;
			sig_dout <= data_mem(to_integer(unsigned(end1))) & data_mem(to_integer(unsigned(end1)+1)) & 
					data_mem(to_integer(unsigned(end1)+2)) & data_mem(to_integer(unsigned(end1)+3));
		else
			sig_dout <= (others => '0');
		end if;
	end process;
	
	dout <= sig_dout;
	
end arch_cache_instrucoes;